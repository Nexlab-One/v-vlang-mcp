module tools

import json
import mcp
import server

// Tool registry maps method names to handler functions
pub type ToolHandler = fn (params mcp.JsonAny, mut docs_server server.VDocumentationServer) string

pub struct ToolRegistry {
mut:
	handlers map[string]ToolHandler
}

pub fn new_tool_registry() ToolRegistry {
	mut registry := ToolRegistry{
		handlers: map[string]ToolHandler{}
	}
	registry.register_all()
	return registry
}

fn (mut r ToolRegistry) register_all() {
	r.handlers['get_v_documentation'] = handle_get_v_documentation
	r.handlers['search_v_docs'] = handle_search_v_docs
	r.handlers['list_v_examples'] = handle_list_v_examples
	r.handlers['get_v_example'] = handle_get_v_example
	r.handlers['search_v_examples'] = handle_search_v_examples
	r.handlers['list_v_stdlib_modules'] = handle_list_v_stdlib_modules
	r.handlers['get_v_module_info'] = handle_get_v_module_info
	r.handlers['explain_v_syntax'] = handle_explain_v_syntax
	r.handlers['get_v_quick_reference'] = handle_get_v_quick_reference
	r.handlers['get_v_config'] = handle_get_v_config
	r.handlers['clear_v_cache'] = handle_clear_v_cache
	r.handlers['list_v_ui_examples'] = handle_list_v_ui_examples
	r.handlers['get_v_ui_example'] = handle_get_v_ui_example
	r.handlers['search_v_ui_examples'] = handle_search_v_ui_examples
	r.handlers['get_v_help'] = handle_get_v_help
}

pub fn (r &ToolRegistry) call_tool(method string, params mcp.JsonAny, mut docs_server server.VDocumentationServer) !string {
	handler := r.handlers[method] or {
		return error('Method not found: ${method}')
	}
	return handler(params, mut docs_server)
}

// Tool handlers

fn handle_get_v_documentation(params mcp.JsonAny, mut docs_server server.VDocumentationServer) string {
	if !docs_server.path_status.docs {
		return '# V Documentation - Not Available\n\nDocumentation is not available. Check V_REPO_PATH environment variable.'
	}

	section_param := mcp.extract_optional_string_param(params, 'section')
	
	sections_json := docs_server.get_documentation_sections()
	sections := json.decode(map[string]string, sections_json) or {
		return '# V Documentation - Error\n\nFailed to parse documentation sections.'
	}

	if 'error' in sections {
		return '# V Documentation - Error\n\n${sections['error']}'
	}

	if section := section_param {
		if section in sections {
			section_content := sections[section] or { '' }
			return '# ${section}\n\n${section_content}'
		} else {
		mut available := []string{}
		keys := sections.keys()
		for key in keys {
			available << key
		}
		return '# Section Not Found\n\nSection "${section}" not found. Available sections: ${available.join(', ')}'
		}
	}

	// Return overview
	mut output := '# V Programming Language Documentation\n\n'
	output += 'Documentation loaded successfully (${sections.len} sections available)\n\n'
	output += '**Available sections:**\n\n'
	for sec in sections.keys() {
		output += '- ${sec}\n'
	}
	output += '\n**Usage:** `get_v_documentation(section_name)` to get specific sections.'
	return output
}

fn handle_search_v_docs(params mcp.JsonAny, mut docs_server server.VDocumentationServer) string {
	query_param := mcp.extract_string_param(params, 'query') or {
		return 'Error: Query parameter is required'
	}

	results_json := docs_server.search_documentation(query_param)
	results := json.decode([]map[string]mcp.JsonAny, results_json) or {
		return 'Error: Failed to parse search results'
	}

	if results.len == 0 {
		return 'No results found for "${query_param}" in V documentation.'
	}

	mut output := '# Search Results for "${query_param}"\n\n'
	mut successful_results := []map[string]mcp.JsonAny{}
	for r in results {
		if 'error' !in r {
			successful_results << r
		}
	}

	if successful_results.len > 0 {
		output += 'Found ${successful_results.len} matches (showing top 10):\n\n'
		max_show := if successful_results.len > 10 { 10 } else { successful_results.len }
		for i := 0; i < max_show; i++ {
			result := successful_results[i].clone()
			file_val := match result['file'] {
				string { result['file'] as string }
				else { 'unknown' }
			}
			line_val := match result['line'] {
				mcp.JsonAnyInt { int(result['line'] as mcp.JsonAnyInt) }
				else { 0 }
			}
			content_val := match result['content'] {
				string { result['content'] as string }
				else { '' }
			}
			context_val := match result['context'] {
				string { result['context'] as string }
				else { '' }
			}
			output += '**File:** ${file_val}\n'
			output += '**Line ${line_val}:** ${content_val}\n'
			output += '**Context:**\n```\n${context_val}\n```\n\n'
		}
	} else {
		for r in results {
			if 'error' in r {
				error_val := match r['error'] {
					string { r['error'] as string }
					else { 'Unknown error' }
				}
				output += 'Error: ${error_val}\n\n'
			}
		}
	}

	return output
}

fn handle_list_v_examples(params mcp.JsonAny, mut docs_server server.VDocumentationServer) string {
	if !docs_server.path_status.examples {
		return '# V Examples - Not Available\n\nExamples directory not found. Check V_REPO_PATH environment variable.'
	}

	examples_json := docs_server.get_examples_list()
	examples := json.decode([]map[string]string, examples_json) or {
		return '# Examples Error\n\nFailed to parse examples list.'
	}

	if examples.len == 0 {
		return '# No Examples Found\n\nNo V examples were found.'
	}

	mut valid_examples := []map[string]string{}
	for ex in examples {
		if 'error' !in ex {
			valid_examples << ex
		}
	}

	mut output := '# V Programming Examples\n\n'
	if valid_examples.len > 0 {
		output += 'Found ${valid_examples.len} examples\n\n'
		max_show := if valid_examples.len > 20 { 20 } else { valid_examples.len }
		for i := 0; i < max_show; i++ {
			ex := valid_examples[i].clone()
			output += '**${ex['name']}**\n'
			output += '- Path: ${ex['path']}\n'
			output += '- Description: ${ex['description']}\n\n'
		}
		if valid_examples.len > 20 {
			output += '\n*Showing first 20 of ${valid_examples.len} examples.*\n'
		}
		output += '*Use `get_v_example(name)` to see the full code for any example.*'
	} else {
		output += 'No valid examples could be loaded.'
	}

	return output
}

fn handle_get_v_example(params mcp.JsonAny, mut docs_server server.VDocumentationServer) string {
	example_name_param := mcp.extract_string_param(params, 'example_name') or {
		return 'Error: example_name parameter is required'
	}

	result_json := docs_server.get_example_content(example_name_param)
	result := json.decode(map[string]string, result_json) or {
		return 'Error: Failed to parse example result'
	}

	if 'error' in result {
		return '# Example Not Found\n\nExample "${example_name_param}" not found.\n\nError: ${result['error']}\n\nUse `list_v_examples()` to see all available examples.'
	}

	mut output := '# V Example: ${result['name']}\n\n'
	output += '**Path:** ${result['path']}\n\n'
	output += '## Source Code\n\n'
	output += '```v\n${result['content']}\n```\n'

	return output
}

fn handle_search_v_examples(params mcp.JsonAny, mut docs_server server.VDocumentationServer) string {
	query_param := mcp.extract_string_param(params, 'query') or {
		return 'Error: Query parameter is required'
	}

	results_json := docs_server.search_examples(query_param)
	results := json.decode([]map[string]mcp.JsonAny, results_json) or {
		return 'Error: Failed to parse search results'
	}

	if results.len == 0 {
		return 'No examples found containing "${query_param}".'
	}

	mut output := '# Examples containing "${query_param}"\n\n'
	mut successful_results := []map[string]mcp.JsonAny{}
	for r in results {
		if 'error' !in r {
			successful_results << r
		}
	}

	if successful_results.len > 0 {
		output += 'Found ${successful_results.len} matches across examples:\n\n'
		max_show := if successful_results.len > 15 { 15 } else { successful_results.len }
		for i := 0; i < max_show; i++ {
			result := successful_results[i].clone()
			file_val := match result['file'] {
				string { result['file'] as string }
				else { 'unknown' }
			}
			line_val := match result['line'] {
				mcp.JsonAnyInt { int(result['line'] as mcp.JsonAnyInt) }
				else { 0 }
			}
			content_val := match result['content'] {
				string { result['content'] as string }
				else { '' }
			}
			output += '**File:** ${file_val}\n'
			output += '**Line ${line_val}:** ${content_val}\n\n'
		}
	}

	return output
}

fn handle_list_v_stdlib_modules(params mcp.JsonAny, mut docs_server server.VDocumentationServer) string {
	modules_json := docs_server.get_stdlib_modules()
	modules := json.decode([]map[string]string, modules_json) or {
		return 'Error: Failed to parse modules list'
	}

	if modules.len == 0 {
		return 'No standard library modules found.'
	}

	mut output := '# V Standard Library Modules\n\n'
	for mod in modules {
		if 'error' !in mod {
			output += '**${mod['name']}**\n'
			output += '- Description: ${mod['description']}\n\n'
		}
	}

	output += '\nUse `get_v_module_info(module_name)` to get detailed information about a specific module.'
	return output
}

fn handle_get_v_module_info(params mcp.JsonAny, mut docs_server server.VDocumentationServer) string {
	module_name_param := mcp.extract_string_param(params, 'module_name') or {
		return 'Error: module_name parameter is required'
	}

	result_json := docs_server.get_module_info(module_name_param)
	result := json.decode(map[string]mcp.JsonAny, result_json) or {
		return 'Error: Failed to parse module info'
	}

	if 'error' in result {
		error_val := match result['error'] {
			string { result['error'] as string }
			else { 'Unknown error' }
		}
		return 'Error: ${error_val}\n\nUse `list_v_stdlib_modules()` to see available modules.'
	}

	mut output := '# V Standard Library Module: ${module_name_param}\n\n'

	if 'readme' in result {
		readme_val := match result['readme'] {
			string { result['readme'] as string }
			else { '' }
		}
		if readme_val != '' {
			output += '## Documentation\n\n'
			output += readme_val
			output += '\n\n'
		}
	}

	if 'files' in result {
		files_val := match result['files'] {
			[]mcp.JsonAny { result['files'] as []mcp.JsonAny }
			else { []mcp.JsonAny{} }
		}
		if files_val.len > 0 {
			output += '## Files\n\n'
			max_show := if files_val.len > 10 { 10 } else { files_val.len }
			for i := 0; i < max_show; i++ {
				file_info := match files_val[i] {
					map[string]mcp.JsonAny { files_val[i] as map[string]mcp.JsonAny }
					else { map[string]mcp.JsonAny{} }
				}
				name_val := match file_info['name'] {
					string { file_info['name'] as string }
					else { 'unknown' }
				}
				size_val := match file_info['size'] {
					mcp.JsonAnyInt { int(file_info['size'] as mcp.JsonAnyInt) }
					else { 0 }
				}
				path_val := match file_info['path'] {
					string { file_info['path'] as string }
					else { 'unknown' }
				}
				output += '- **${name_val}** (${size_val} bytes)\n'
				output += '  - Path: ${path_val}\n'
			}
			if files_val.len > 10 {
				output += '\n*... and ${files_val.len - 10} more files*\n'
			}
		}
	}

	return output
}

fn handle_explain_v_syntax(params mcp.JsonAny, mut docs_server server.VDocumentationServer) string {
	feature_param := mcp.extract_string_param(params, 'feature') or {
		return 'Error: feature parameter is required'
	}

	feature := feature_param.to_lower().trim_space()
	
	features := get_v_syntax_features()
	
	if feature in features {
		return features[feature]
	}

	mut available := []string{}
	keys := features.keys()
	for key in keys {
		available << key
	}
	return 'Feature "${feature_param}" not found. Available features: ${available.join(', ')}\n\nUse `search_v_docs("${feature_param}")` to search documentation for this topic.'
}

fn handle_get_v_quick_reference(params mcp.JsonAny, mut docs_server server.VDocumentationServer) string {
	return get_v_quick_reference_content()
}

fn handle_get_v_config(params mcp.JsonAny, mut docs_server server.VDocumentationServer) string {
	stats := docs_server.get_cache_stats()
	
	mut output := '# V MCP Server Configuration\n\n'
	output += '**V Repository Path:** ${docs_server.config.v_repo_path}\n'
	if docs_server.config.v_ui_path != '' {
		output += '**V UI Path:** ${docs_server.config.v_ui_path}\n'
	} else {
		output += '**V UI Path:** Not configured\n'
	}
	output += '**Cache TTL:** ${docs_server.config.cache_ttl_seconds}s\n'
	output += '**Max Search Results:** ${docs_server.config.max_search_results}\n'
	output += '**Log Level:** ${docs_server.config.log_level}\n\n'
	output += '**Path Status:**\n'
	output += '- Documentation: ${if docs_server.path_status.docs { 'Available' } else { 'Not available' }}\n'
	output += '- Examples: ${if docs_server.path_status.examples { 'Available' } else { 'Not available' }}\n'
	output += '- Standard Library: ${if docs_server.path_status.stdlib { 'Available' } else { 'Not available' }}\n'
	output += '- V UI: ${if docs_server.path_status.v_ui { 'Available' } else { 'Not available' }}\n'
	output += '- V UI Examples: ${if docs_server.path_status.v_ui_examples { 'Available' } else { 'Not available' }}\n\n'
	output += '**Cache Statistics:**\n'
	output += '- Current cache entries: ${stats['entries']}\n'
	output += '- Cache TTL: ${stats['ttl_seconds']}s\n'

	return output
}

fn handle_clear_v_cache(params mcp.JsonAny, mut docs_server server.VDocumentationServer) string {
	result_json := docs_server.clear_cache()
	result := json.decode(map[string]int, result_json) or {
		return 'Error: Failed to parse cache clear result'
	}

	mut output := '# Cache Cleared\n\n'
	output += 'Cleared ${result['cleared_entries']} cache entries\n\n'
	output += '**Statistics:**\n'
	output += '- Cache entries cleared: ${result['cleared_entries']}\n'
	output += '- Timestamp entries cleared: ${result['cleared_timestamps']}\n\n'
	output += 'Next requests will reload content from the V repository.'

	return output
}

fn handle_list_v_ui_examples(params mcp.JsonAny, mut docs_server server.VDocumentationServer) string {
	if !docs_server.path_status.v_ui_examples {
		return json.encode({
			'error': 'V UI examples are not available'
			'message': 'V UI repository not found or examples directory missing. Make sure the v-ui submodule is initialized.'
		})
	}

	examples_json := docs_server.get_v_ui_examples_list()
	return examples_json
}

fn handle_get_v_ui_example(params mcp.JsonAny, mut docs_server server.VDocumentationServer) string {
	example_name_param := mcp.extract_string_param(params, 'example_name') or {
		return json.encode({
			'error': 'example_name parameter is required'
		})
	}

	if !docs_server.path_status.v_ui_examples {
		return json.encode({
			'error': 'V UI examples are not available'
			'message': 'V UI repository not found or examples directory missing.'
		})
	}

	return docs_server.get_v_ui_example_content(example_name_param)
}

fn handle_search_v_ui_examples(params mcp.JsonAny, mut docs_server server.VDocumentationServer) string {
	query_param := mcp.extract_string_param(params, 'query') or {
		return json.encode({
			'error': 'Query parameter is required'
		})
	}

	if !docs_server.path_status.v_ui_examples {
		return json.encode({
			'error': 'V UI examples are not available'
			'message': 'V UI repository not found or examples directory missing.'
		})
	}

	vui_search_results_json := docs_server.search_v_ui_examples(query_param)
	vui_search_results := json.decode([]map[string]mcp.JsonAny, vui_search_results_json) or {
		return json.encode({
			'error': 'Failed to parse search results'
		})
	}

	// Return result as map with mixed types - encode manually
	mut vui_result_map := map[string]mcp.JsonAny{}
	vui_result_map['query'] = mcp.JsonAny(query_param)
	vui_result_map['count'] = mcp.JsonAny(mcp.JsonAnyInt(vui_search_results.len))
	mut vui_results_array := []mcp.JsonAny{}
		for r in vui_search_results {
			vui_results_array << r
		}
	vui_result_map['results'] = mcp.JsonAny(vui_results_array)
	return json.encode(vui_result_map)
}

fn handle_get_v_help(params mcp.JsonAny, mut docs_server server.VDocumentationServer) string {
	return get_v_help_content()
}

// Helper functions for static content

fn get_v_syntax_features() map[string]string {
	return {
		'variables': '# V Variables\n\nV supports several types of variables:\n\n## Declaration and Initialization\n```v\nname := \'Bob\'  // Inferred type string\nage := 20       // Inferred type int\nis_adult := true // Inferred type bool\n```\n\n## Explicit Type Declaration\n```v\nmut name string = \'Bob\'  // Mutable variable\nage int = 20            // Immutable variable\n```\n\n## Constants\n```v\nconst pi = 3.14159\nconst (\n    rate = 0.05\n    days = 365\n)\n```\n'
		'arrays': '# V Arrays\n\n## Declaration and Initialization\n```v\nmut numbers := [1, 2, 3]     // Inferred type []int\nnames := [\'Alice\', \'Bob\']    // []string\nempty := []int{}             // Empty array\n```\n\n## Array Operations\n```v\nnumbers << 4                 // Append element\nnumbers << [5, 6]            // Append array\nfirst := numbers[0]          // Access element\nnumbers[1] = 10              // Modify element\nlen := numbers.len           // Get length\n```\n\n## Array Methods\n```v\nnumbers.insert(0, 0)         // Insert at index\nnumbers.delete(1)            // Delete element\nnumbers.reverse()            // Reverse array\nnumbers.sort()               // Sort array\n```\n'
		'structs': r"# V Structs

## Definition
```v
struct User {
    id   int
    name string
    age  int
mut:
    email string  // Mutable field
pub:
    active bool   // Public field
}
```

## Usage
```v
user := User{
    id: 1
    name: 'Alice'
    age: 30
    email: 'alice@example.com'
    active: true
}

// Access fields
println(user.name)    // Alice
user.email = 'new@example.com'  // Modify mutable field
```

## Methods
```v
fn (u User) full_name() string {
    return u.name + ' (ID: ' + u.id.str() + ')'
}

fn (mut u User) deactivate() {
    u.active = false
}
```
"
		'functions': '# V Functions\n\n## Basic Function\n```v\nfn greet(name string) string {\n    return \'Hello, \' + name + \'!\'\n}\n\nmessage := greet(\'World\')\n```\n\n## Multiple Return Values\n```v\nfn divide(a int, b int) (int, int) {\n    quotient := a / b\n    remainder := a % b\n    return quotient, remainder\n}\n\nq, r := divide(10, 3)\n```\n\n## Variadic Functions\n```v\nfn sum(numbers ...int) int {\n    mut total := 0\n    for num in numbers {\n        total += num\n    }\n    return total\n}\n\nresult := sum(1, 2, 3, 4, 5)\n```\n'
		'control_flow': '# V Control Flow\n\n## If Statements\n```v\nage := 18\nif age >= 18 {\n    println(\'Adult\')\n} else if age >= 13 {\n    println(\'Teenager\')\n} else {\n    println(\'Child\')\n}\n```\n\n## If as Expression\n```v\nmax := if a > b { a } else { b }\nstatus := if user.active { \'Active\' } else { \'Inactive\' }\n```\n\n## Match Statement\n```v\ncolor := \'red\'\nmatch color {\n    \'red\' { println(\'Stop!\') }\n    \'yellow\' { println(\'Caution!\') }\n    \'green\' { println(\'Go!\') }\n    else { println(\'Unknown color\') }\n}\n```\n\n## For Loops\n```v\n// Basic loop\nfor i in 0..10 {\n    println(i)\n}\n\n// Loop over array\nfruits := [\'apple\', \'banana\', \'cherry\']\nfor fruit in fruits {\n    println(fruit)\n}\n\n// Loop with index\nfor i, fruit in fruits {\n    println(i.str() + \': \' + fruit)\n}\n```\n'
		'modules': '# V Modules\n\n## Module Declaration\nEach V file belongs to a module. The module name is the same as the folder name.\n\n## Importing Modules\n```v\nimport os\nimport utils.math\nimport utils.string as str_utils\n```\n\n## Selective Imports\n```v\nimport os { read_file, write_file }\nimport utils.math { add, multiply as mul }\n```\n'
		'error_handling': '# V Error Handling\n\n## Option Types\n```v\nfn find_user(id int) ?User {\n    if id < 0 {\n        return none\n    }\n    return User{ id: id, name: \'User \' + id.str() }\n}\n\n// Usage\nuser := find_user(123) or {\n    println(\'User not found\')\n    return\n}\nprintln(user.name)\n```\n\n## Error Types\n```v\nfn risky_operation() !string {\n    if rand.intn(2) == 0 {\n        return error(\'Something went wrong\')\n    }\n    return \'Success!\'\n}\n\n// Usage\nresult := risky_operation() or {\n    println(\'Error: \' + err.str())\n    exit(1)\n}\nprintln(result)\n```\n'
		'concurrency': '# V Concurrency\n\n## Goroutines\n```v\nfn worker(id int) {\n    println(\'Worker \' + id.str() + \' starting\')\n    time.sleep(1 * time.second)\n    println(\'Worker \' + id.str() + \' done\')\n}\n\nfn main() {\n    for i in 1..5 {\n        go worker(i)\n    }\n    time.sleep(2 * time.second)\n}\n```\n\n## Channels\n```v\nfn producer(ch chan int) {\n    for i in 1..10 {\n        ch <- i\n        time.sleep(100 * time.millisecond)\n    }\n    ch.close()\n}\n\nfn consumer(ch chan int) {\n    for {\n        if val := <-ch {\n            println(\'Received: \' + val.str())\n        } else {\n            break  // Channel closed\n        }\n    }\n}\n\nfn main() {\n    ch := chan int{}\n    go producer(ch)\n    consumer(ch)\n}\n```\n'
	}
}

fn get_v_quick_reference_content() string {
	return '# V Programming Language Quick Reference\n\n## Basic Syntax\n```v\n// Hello World\nfn main() {\n    println(\'Hello, World!\')\n}\n\n// Variables\nname := \'Bob\'  // Inferred type\nage int = 20   // Explicit type\nmut count := 0 // Mutable\n\n// Arrays\nnumbers := [1, 2, 3]\nnumbers << 4  // Append\nfirst := numbers[0]\n\n// Structs\nstruct User {\n    id   int\n    name string\n}\n\nuser := User{ id: 1, name: \'Alice\' }\n\n// Functions\nfn greet(name string) string {\n    return \'Hello, \' + name + \'!\'\n}\n\n// Control Flow\nif age >= 18 {\n    println(\'Adult\')\n}\n\nfor i in 0..10 {\n    println(i)\n}\n\n// Error Handling\nresult := risky_op() or {\n    println(\'Error: \' + err.str())\n    return\n}\n\n// Concurrency\ngo worker()\nch := chan int{}\nch <- 42\nvalue := <-ch\n```\n\nFor more detailed information, use the other tools available.'
}

fn get_v_help_content() string {
	return '# V MCP Server Help\n\nThe V MCP Server provides comprehensive access to V programming language resources.\n\n## Available Tools\n\n### Documentation Tools\n- **`get_v_documentation([section])`** - Get V documentation, optionally for a specific section\n- **`search_v_docs(query)`** - Search through V documentation\n\n### Code Examples\n- **`list_v_examples()`** - List all available V code examples\n- **`get_v_example(name)`** - Get complete source code for a specific example\n- **`search_v_examples(query)`** - Search through example code\n\n### Standard Library\n- **`list_v_stdlib_modules()`** - List all V standard library modules\n- **`get_v_module_info(module_name)`** - Get detailed info about a specific module\n\n### V UI Examples\n- **`list_v_ui_examples()`** - List all available V UI code examples\n- **`get_v_ui_example(name)`** - Get complete source code for a specific V UI example\n- **`search_v_ui_examples(query)`** - Search through V UI example code\n\n### Language Reference\n- **`explain_v_syntax(feature)`** - Explain V language features\n- **`get_v_quick_reference()`** - Get quick V syntax reference\n\n### Configuration & Cache\n- **`get_v_config()`** - Show current server configuration and cache statistics\n- **`clear_v_cache()`** - Clear cached content for fresh results\n\n### Help & Discovery\n- **`get_v_help()`** - Show this help information\n\n## Usage Tips\n\n1. Start with the basics: Use `get_v_quick_reference()` to learn essential syntax\n2. Explore examples: Use `list_v_examples()` to see practical code\n3. Search documentation: Use `search_v_docs()` for specific topics\n4. Learn features: Use `explain_v_syntax()` for detailed explanations\n5. Browse stdlib: Use `list_v_stdlib_modules()` to explore available modules\n6. Check configuration: Use `get_v_config()` to verify server settings\n7. Clear cache when needed: Use `clear_v_cache()` after V repository updates'
}
